LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY deco IS
	PORT(DEC: IN INTEGER RANGE 0 TO 9; -- ENTRADA ENTRE EL 0 Y 9
	SEG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)); -- DISPLAY 7 SEG
END deco;

ARCHITECTURE BEAS OF deco IS
BEGIN
	-- Decodificador de decimal a 7 seg
	WITH DEC SELECT
		SEG <= 	"00000011" WHEN 0, -- 0
					"10011111" WHEN 1, -- 1
					"00100101" WHEN 2, -- 2
					"00001101" WHEN 3, -- 3
					"10011001" WHEN 4, -- 4
					"01001001" WHEN 5, -- 5
					"01000001" WHEN 6, -- 6
					"00011111" WHEN 7, -- 7
					"00000001" WHEN 8, -- 8
					"00001001" WHEN 9, -- 9
					"11111111" WHEN OTHERS; -- OTROS CASOS

END BEAS;