LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;

ENTITY decop IS
	PORT(DEC: IN INTEGER RANGE 0 TO 9; -- ENTRADA ENTRE EL 0 Y 9
	SEG: OUT STD_LOGIC_VECTOR(7 DOWNTO 0)); -- DISPLAY 7 SEG
END decop;

ARCHITECTURE BEAS OF decop IS
BEGIN
	-- Decodificador de decimal a 7 seg
	WITH DEC SELECT
		SEG <= 	"00000010" WHEN 0, -- 0
					"10011110" WHEN 1, -- 1
					"00100100" WHEN 2, -- 2
					"00001100" WHEN 3, -- 3
					"10011000" WHEN 4, -- 4
					"01001000" WHEN 5, -- 5
					"01000000" WHEN 6, -- 6
					"00011110" WHEN 7, -- 7
					"00000000" WHEN 8, -- 8
					"00001000" WHEN 9, -- 9
					"11111110" WHEN OTHERS; -- OTROS CASOS

END BEAS;